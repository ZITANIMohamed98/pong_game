//=============================================================================================
//    Main contributors
//      - Adam Luczak         <mailto:aluczak@multimedia.edu.pl>
//=============================================================================================
`default_nettype none
//---------------------------------------------------------------------------------------------
`timescale 1ns / 1ns                            
//=============================================================================================
module dev_i2c_phy_bit
(
input  wire	        clk,
input  wire	        tick,
input  wire         rst,   

input  wire         i_stb,
input  wire         i_dir,
input  wire  [1:0]  i_bit,
output wire         i_ack,
output wire         i_rdy,

output wire         o_val,
output wire         o_lde,
output wire         o_bit,

// I2C bus
inout  wire         i2c_sda,
output wire         i2c_scl
);
//==============================================================================================
// local param
//==============================================================================================
//==============================================================================================
// variables
//==============================================================================================   
reg   [1:0] bit_data;      
reg   [1:0] bit_phase;
reg         bit_dir;
reg         bit_run;
reg         bit_rdy;
//---------------------------------------------------------------------------------------------- 
reg         sda_0; 
reg         sen_0; 
reg         scl_0; 
//---------------------------------------------------------------------------------------------- 
reg         sda_1; 
reg         sen_1; 
reg         scl_1; 
//---------------------------------------------------------------------------------------------- 
reg         sda_2; 
//---------------------------------------------------------------------------------------------- 
reg         sda_3;         
reg         val_3;
reg         lde_3;
//==============================================================================================
// control flags
//==============================================================================================
wire          f_ld_start                =                             i_stb & i_bit    == 2'b10;
wire          f_ld_bit                  =                             i_stb & i_bit[1] == 1'b0;
wire          f_ld_stop                 =                             i_stb & i_bit    == 2'b11;
//---------------------------------------------------------------------------------------------- 
wire          f_lde                     =                                         i_stb && tick;
wire          f_inc                     =                              bit_phase!=2'b11 && tick;
wire          f_rdy                     =                              bit_phase==2'b11;
wire          f_clr                     =                              bit_phase==2'b11 && tick;
//---------------------------------------------------------------------------------------------- 
wire          f_sample                  =                              bit_phase==2'b01 && tick;
wire          f_out_tick                =                              bit_phase==2'b10 && tick;
//==============================================================================================
// BIT SENDER
//==============================================================================================
always@(posedge clk or posedge rst)
  if(rst)                   bit_data    <=                                                2'b11;
  else if(f_lde)            bit_data    <=                                                i_bit;
//---------------------------------------------------------------------------------------------- 
always@(posedge clk or posedge rst)
  if(rst)                   bit_dir     <=                                                 1'b1;
  else if(f_lde)            bit_dir     <=                                                i_dir;
//---------------------------------------------------------------------------------------------- 
always@(posedge clk or posedge rst)
  if(rst)                   bit_run     <=                                                 1'b0;
  else if(f_lde)            bit_run     <=                                                 1'b1;
  else if(f_clr)            bit_run     <=                                                 1'b0;
//---------------------------------------------------------------------------------------------- 
always@(posedge clk or posedge rst)
  if(rst)                   bit_phase   <=                                                2'b11;
  else if(f_lde)            bit_phase   <=                                                2'b00;
  else if(f_inc)            bit_phase   <=                                     bit_phase + 2'd1;
//----------------------------------------------------------------------------------------------       
always@(posedge clk or posedge rst)
  if(rst)                   bit_rdy     <=                                                 1'b1;
  else if(f_lde)            bit_rdy     <=                                                 1'b0;
  else if(f_rdy)            bit_rdy     <=                                                 1'b1;
//---------------------------------------------------------------------------------------------- 
assign                      i_ack        =                                                f_lde;
assign                      i_rdy        =                                              bit_rdy;
//----------------------------------------------------------------------------------------------       
// i2c clk waveform
//---------------------------------------------------------------------------------------------- 
always@(posedge clk or posedge rst)
  if(rst)                   scl_0       <=                                                 1'b1;   
  else if(bit_data==2'b00 && bit_run) // bit 0 
    case(bit_phase)
    2'd0 :                  scl_0       <=                                                 1'b0;
    2'd1 :                  scl_0       <=                                                 1'b1;
    2'd2 :                  scl_0       <=                                                 1'b1;
    2'd3 :                  scl_0       <=                                                 1'b0;
    endcase 
  else if(bit_data==2'b01 && bit_run) // bit 1 
    case(bit_phase)
    2'd0 :                  scl_0       <=                                                 1'b0;
    2'd1 :                  scl_0       <=                                                 1'b1;
    2'd2 :                  scl_0       <=                                                 1'b1;
    2'd3 :                  scl_0       <=                                                 1'b0;
    endcase 
  else if(bit_data==2'b10 && bit_run) // start bit 
    case(bit_phase)
    2'd0 :                  scl_0       <=                                                 1'b1;
    2'd1 :                  scl_0       <=                                                 1'b1;
    2'd2 :                  scl_0       <=                                                 1'b1;
    2'd3 :                  scl_0       <=                                                 1'b0;
    endcase 
  else if(bit_data==2'b11 && bit_run) // stop bit 
    case(bit_phase)
    2'd0 :                  scl_0       <=                                                 1'b0;
    2'd1 :                  scl_0       <=                                                 1'b1;
    2'd2 :                  scl_0       <=                                                 1'b1;
    2'd3 :                  scl_0       <=                                                 1'b1;
    endcase 
  else                      scl_0       <=                                                scl_0;                
//---------------------------------------------------------------------------------------------- 
// i2c data waveform
//---------------------------------------------------------------------------------------------- 
always@(posedge clk or posedge rst)
  if(rst)                   sda_0       <=                                                 1'b1;   
  else if(bit_data==2'b00 && bit_run) // bit 0
    case(bit_phase)
    2'd0 :                  sda_0       <=                                                 1'b0;
    2'd1 :                  sda_0       <=                                                 1'b0;
    2'd2 :                  sda_0       <=                                                 1'b0;
    2'd3 :                  sda_0       <=                                                 1'b0;
    endcase 
  else if(bit_data==2'b01 && bit_run) // bit 1
    case(bit_phase)
    2'd0 :                  sda_0       <=                                                 1'b1;
    2'd1 :                  sda_0       <=                                                 1'b1;
    2'd2 :                  sda_0       <=                                                 1'b1;
    2'd3 :                  sda_0       <=                                                 1'b1;
    endcase 
  else if(bit_data==2'b10 && bit_run) // start bit 
    case(bit_phase)
    2'd0 :                  sda_0       <=                                                 1'b1;
    2'd1 :                  sda_0       <=                                                 1'b1;
    2'd2 :                  sda_0       <=                                                 1'b0;
    2'd3 :                  sda_0       <=                                                 1'b0;
    endcase 
  else if(bit_data==2'b11 && bit_run) // stop bit 
    case(bit_phase)
    2'd0 :                  sda_0       <=                                                 1'b0;
    2'd1 :                  sda_0       <=                                                 1'b0;
    2'd2 :                  sda_0       <=                                                 1'b1;
    2'd3 :                  sda_0       <=                                                 1'b1;
    endcase 
  else                      sda_0       <=                                                scl_0;                
//----------------------------------------------------------------------------------------------                       
// tristate line SDA "enabled" signal                                                                                  
//---------------------------------------------------------------------------------------------- 
always@(posedge clk or posedge rst)
  if(rst)                   sen_0       <=                                                 1'b1;
  else                      sen_0       <=                                              bit_dir;    
//==============================================================================================
// I/O buffer 
//==============================================================================================
always@(posedge clk or posedge rst)
  if(rst)                   scl_1        <=                                               1'b1;
  else                      scl_1        <=                                               scl_0;
//---------------------------------------------------------------------------------------------- 
always@(posedge clk or posedge rst)
  if(rst)                   sda_1        <=                                               1'b1;
  else                      sda_1        <=                                               sda_0;
//---------------------------------------------------------------------------------------------- 
always@(posedge clk or posedge rst)
  if(rst)                   sen_1        <=                                               1'b1;
  else                      sen_1        <=                                               sen_0;
//==============================================================================================
// i2c output
//==============================================================================================
assign                    i2c_sda         = (sen_1==1'b0) ?                        1'bz : sda_1;
assign                    i2c_scl         =                                               scl_1;
//==============================================================================================
// input I/O
//==============================================================================================
always@(posedge clk)        sda_2        <=                                             i2c_sda;
//---------------------------------------------------------------------------------------------- 
// input bit sampling
//---------------------------------------------------------------------------------------------- 
always@(posedge clk or posedge rst)                                                                         
  if(rst)                   sda_3        <=                                                1'b1;                                                          
  else if(f_sample)         sda_3        <=                                               sda_2;
//---------------------------------------------------------------------------------------------- 
always@(posedge clk or posedge rst)
  if(rst)                   val_3        <=                                                1'b0;
  else if(f_sample)         val_3        <=                                                1'b1;
  else if(f_lde)            val_3        <=                                                1'b0;
//---------------------------------------------------------------------------------------------- 
always@(posedge clk or posedge rst)                                                                         
  if(rst)                   lde_3        <=                                                1'b0;
  else if(f_out_tick)       lde_3        <=                                                1'b1;
  else                      lde_3        <=                                                1'b0;
//==============================================================================================
// output
//==============================================================================================
assign                      o_val        =                                                val_3;
assign                      o_lde        =                                                lde_3;
assign                      o_bit        =                                                sda_3;
//==============================================================================================
endmodule









